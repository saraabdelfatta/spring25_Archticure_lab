`timescale 1ns / 1ps



module inv(
input x,
output y
    );
    
    assign y = ~x;
endmodule
